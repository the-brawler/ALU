module testbench_ALU();
    reg [31:0] A, B;
	reg [3:0] Operator;
	reg [5:0] n;
    wire [31:0] Result;
 
    alu U1 (.A(A),.B(B),.Operator(Operator),.n(n),.Result(Result));
    
    initial
	begin

		A = 32'b01100111000010000101000110000110;
		B = 32'b01010101101101111101010011000111;
		n=6'd32;
		Operator=4'b0000;
		#100
					  
			 
		A = 32'b10111110001010111011010011111100;
		B = 32'b00011011000000001100100110100001;
		n=6'd3;
		Operator=4'b0001;
		#100 
					  
			 
		A = 32'b10011101111100111011011000111001;
		B = 32'b01010000111001001001110000010100;
		n=6'd0;
		Operator=4'b0010;
		#100 
			 
		A = 32'b00100001101110001001100011010101;
		B = 32'b10101000100111110111101001011101;
		n=6'd1;
		Operator=4'b0011;
		#100 
					  
			 
		A = 32'b00110101101110110010000111000100;
		B = 32'b10001011010100000001100000110111;
		n=6'd4;
		Operator=4'b0100;
		#100 
					  
			 
		A = 32'b10001011100111001011101111010101;
		B = 32'b10011010010100010001111100000000;
		n=6'd13;
		Operator=4'b0101;
		#100 
					  
			 
		A = 32'b10100101000011101110000101100111;
		B = 32'b10010100111100111110010000001000;
		n=6'd9;
		Operator=4'b0110;
		#100 
					  
			 
		A = 32'b00101011100001011000110011000101;
		B = 32'b11010010010011100000010111100111;
		n=6'd12;
		Operator=4'b0111;
		#100
					  
			 
		A = 32'b10110101100101101100110010100010;
		B = 32'b00000101000111000101000101010110;
		n=6'd9;
		Operator=4'b1000;
		#100
					  
			 
		A = 32'b11110011011100101100111000010010;
		B = 32'b01111010011010100110010001100010;
		n=6'd18;
		Operator=4'b1001;
		#100 
					  
			 
		A = 32'b10000010101101100010100110100101;
		B = 32'b00101001000011110010110100110101;
		n=6'd3;
		Operator=4'b1010;
		#100 
					  
			 
		A = 32'b10101000101010101101100011101001;
		B = 32'b10110010010100100001011011101100;
		n=6'd1;
		Operator=4'b0000;
		#100 
					  
			 
		A = 32'b00010100001101011010101100110111;
		B = 32'b11000011011000011000010100111000;
		n=6'd13;
		Operator=4'b0001;
		#100 
					  
			 
		A = 32'b10010100010010101011111100011000;
		B = 32'b00101101110010100111001010010101;
		n=6'd22;
		Operator=4'b0010;
		#100 
					  
			 
		A = 32'b11101101001100010100010001010001;
		B = 32'b11110101100101101010111111001110;
		n=6'd9;
		Operator=4'b0011;
		#100 
					  
			 
		A = 32'b11100011101110100000001010010111;
		B = 32'b01001101111000110101110000101110;
		n=6'd15;
		Operator=4'b0100;
		#100
					  
			 
		A = 32'b01001010000001100110000111001111;
		B = 32'b01011011100010000110001100010001;
		n=6'd21;
		Operator=4'b0101;
		#100 
					  
			 
		A = 32'b01110000010010111110111110100110;
		B = 32'b11110010000110000111011110110001;
		n=6'd3;
		Operator=4'b0110;
		#100
			 
		A = 32'b00100010101001011010010111101000;
		B = 32'b00010010100100101010110100000100;
		n=6'd4;
        Operator=4'b0111;		
		#100
					  
			 
		A = 32'b10111110100101001001111000100100;
		B = 32'b01011111100010010000001010110000;
		n=6'd16;
		Operator=4'b1000;
		#100
					  
			 
		A = 32'b11011001100110010100110011010011;
		B = 32'b10100111111110100100100000011101;
		n=6'd6;
		Operator=4'b1001;
		#100 
					  
			 
		A = 32'b10111010000100001100101000111110;
		B = 32'b11001011001101010110110010110100;
		n=6'd15;
		Operator=4'b1010;
		#100
					  
			 
		A = 32'b01100110101000001110100111010101;
		B = 32'b10111111001010000100111110101101;
		n=6'd10;
		Operator=4'b0000;
		#100 
					  
			 
		A = 32'b01110011011010001011101101010010;
		B = 32'b01100010111011000000010000011011;
		n=6'd3;
		Operator=4'b0001;
		#100 
			 
		A = 32'b11110000100111101110010110101101;
		B = 32'b11010110111011011010001001110011;
		n=6'd9;
		Operator=4'b0010;
		#100
					  
			 
		A = 32'b10101101101111001111010001101110;
		B = 32'b10001001011001011011110111011000;
		n=6'd26;
		Operator=4'b0011;
		#100 
					  
			 
		A = 32'b11111001111000011110001101100011;
		B = 32'b11101011101000110011100100001011;
		n=6'd9;
		Operator=4'b0100;
		#100 
					  
			 
		A = 32'b00100110010101110001110000000110;
		B = 32'b00010010111100001001110111010011;
		n=6'd2;
		Operator=4'b0101;
		#100 
			 
		A = 32'b01001111110100000010011000111111;
		B = 32'b10100000101011010111001111110100;
		n=6'd3;
		Operator=4'b0110;
		#100 
			 
		A = 32'b01100000011010000001111110001111;
		B = 32'b00101100110100100010111011100001;
		n=6'd6;
		Operator=4'b0111;
		#100 
					  
			 
		A = 32'b00101011101001010001110111011100;
		B = 32'b10101101110000111000100010011111;
		n=6'd5;
		Operator=4'b1000;
		#100 
					  
			 
		A = 32'b11101010110010000111011011001010;
		B = 32'b11001111011101110010110000000010;
		n=6'd2;
		Operator=4'b1001;
		#100 
					  
			 
		A = 32'b01101010011101000001010001100001;
		B = 32'b01100110101010100101011001010001;
		n=6'd4;
		Operator=4'b1010;
		#100 

					  
			 
		A = 32'b00111101010101111101010100101110;
		B = 32'b10101101011100011111001100110011;
		n=6'd8;
		Operator=4'b0000;
		#100 
					  
			 
		A = 32'b01010111111100001000011101010100;
		B = 32'b11100001110101101111100000001110;
		n=6'd12;
		Operator=4'b0001;
		#100 
					  
			 
		A = 32'b11001100010000100111101010000111;
		B = 32'b00101110010011110010100110011000;
		n=6'd7;
		Operator=4'b0010;
		#100
					  
			 
		A = 32'b10010000001011000001001000011010;
		B = 32'b00111001111011011110100000011001;
		n=6'd4;
		Operator=4'b0011;
		#100 
					  
			 
		A = 32'b01001010110010101010001100111000;
		B = 32'b01011101001001111011000111100011;
		n=6'd2;
		Operator=4'b0100;
		#100 
					  
			 
		A = 32'b11011011110100001101000011110001;
		B = 32'b00011101111101001010101011111100;
		n=6'd14;
		Operator=4'b0101;
		#100
					  
			 
		A = 32'b11001110101101101110010000110010;
		B = 32'b11001110110001110110000010000010;
		n=6'd24;
		Operator=4'b0110;
		
					  
			 
	
end 
endmodule